import nyakuo_pkg::*;

module decoder (
  input logic [6:0] opcode_i,
  output logic instruction
);


endmodule